//
// coding convention dudy December 2018
// (c) Technion IIT, Department of Electrical Engineering 2019 
// generating a letter bitmap 



module GameNameLettersBitMap	(	
					input		logic	clk,
					input		logic	resetN,
					input 	logic	[10:0] offsetX,// offset from top left  position 
					input 	logic	[10:0] offsetY,
					input		logic	InsideRectangle, //input that the pixel is within a bracket 
					input 	logic	[5:0] letter, // digit to display
					
					output	logic				drawingRequest, //output that the pixel should be dispalyed 
					output	logic	[7:0]		RGBout
);
// generating a smily bitmap 

parameter  logic	[7:0] digit_color = 8'hff ; //set the color of the digit 


bit [0:19] [0:15] [0:7] letter_bitmap  = {


{8'b	00000000,// no letter
8'b	00000000,
8'b	00000000,
8'b	00000000,
8'b	00000000,
8'b	00000000,
8'b	00000000,
8'b	00000000,
8'b	00000000,
8'b	00000000,
8'b	00000000,
8'b	00000000,
8'b	00000000,
8'b	00000000,
8'b	00000000,
8'b	00000000},

{8'b  00000000,// -- 0 // P
8'b   00000000,// -- 1
8'b   11111100,// -- 2 ******
8'b   01100110,// -- 3  **  **
8'b   01100110,// -- 4  **  **
8'b   01100110,// -- 5  **  **
8'b   01111100,// -- 6  *****
8'b   01100000,// -- 7  **
8'b   01100000,// -- 8  **
8'b   01100000,// -- 9  **
8'b   01100000,// -- a  **
8'b   11110000,// -- b ****
8'b   00000000,// -- c
8'b   00000000,// -- d
8'b   00000000,// -- e
8'b   00000000},// -- f


{8'b	00000000,// -- 0 // R
8'b	00000000,// -- 1
8'b	11111100,// -- 2 ******
8'b	01100110,// -- 3  **  **
8'b	01100110,// -- 4  **  **
8'b	01100110,// -- 5  **  **
8'b	01111100,// -- 6  *****
8'b	01101100,// -- 7  ** **
8'b	01100110,// -- 8  **  **
8'b	01100110,// -- 9  **  **
8'b	01100110,// -- a  **  **
8'b	11100110,// -- b ***  **
8'b	00000000,//-- c
8'b	00000000,// -- d
8'b	00000000,// -- e
8'b	00000000},// -- f

{8'b	00000000,// -- 0 // E
8'b	00000000,// -- 1
8'b	11111110,// -- 2 *******
8'b	01100110,// -- 3  **  **
8'b	01100010,// -- 4  **   *
8'b	01101000,// -- 5  ** *
8'b	01111000,// -- 6  ****
8'b	01101000,// -- 7  ** *
8'b	01100000,// -- 8  **
8'b	01100010,// -- 9  **   *
8'b	01100110,// -- a  **  **
8'b	11111110,// -- b *******
8'b	00000000,// -- c
8'b	00000000,// -- d
8'b	00000000,// -- e
8'b	00000000},// -- f

{8'b	00000000,// -- 0 // S
8'b	00000000,// -- 1
8'b	01111100,// -- 2  *****
8'b	11000110,// -- 3 **   **
8'b	11000110,// -- 4 **   **
8'b	01100000,// -- 5  **
8'b	00111000,// -- 6   ***
8'b	00001100,// -- 7     **
8'b	00000110,// -- 8      **
8'b	11000110,// -- 9 **   **
8'b	11000110,// -- a **   **
8'b	01111100,// -- b  *****
8'b	00000000,// -- c
8'b	00000000,// -- d
8'b	00000000,// -- e
8'b	00000000},// -- f

{8'b	00000000,// -- 0 // A
8'b	00000000,// -- 1
8'b	00010000,// -- 2    *
8'b	00111000,// -- 3   ***
8'b	01101100,// -- 4  ** **
8'b	11000110,// -- 5 **   **
8'b	11000110,// -- 6 **   **
8'b	11111110,// -- 7 *******
8'b	11000110,// -- 8 **   **
8'b	11000110,// -- 9 **   **
8'b	11000110,// -- a **   **
8'b	11000110,// -- b **   **
8'b	00000000,// -- c
8'b	00000000,// -- d
8'b	00000000,// -- e
8'b	00000000},// -- f

{8'b	00000000,// -- 0 // C
8'b	00000000,// -- 1
8'b	00111100,// -- 2   ****
8'b	01100110,// -- 3  **  **
8'b	11000010,// -- 4 **    *
8'b	11000000,// -- 5 **
8'b	11000000,// -- 6 **
8'b	11000000,// -- 7 **
8'b	11000000,// -- 8 **
8'b	11000010,// -- 9 **    *
8'b	01100110,// -- a  **  **
8'b	00111100,// -- b   ****
8'b	00000000,// -- c
8'b	00000000,// -- d
8'b	00000000,// -- e
8'b	00000000},// -- f

{8'b	00000000,// -- 0 // T
8'b	00000000,// -- 1
8'b	11111111,// -- 2 ********
8'b	11011011,// -- 3 ** ** **
8'b	10011001,// -- 4 *  **  *
8'b	00011000,// -- 5    **
8'b	00011000,// -- 6    **
8'b	00011000,// -- 7    **
8'b	00011000,// -- 8    **
8'b	00011000,// -- 9    **
8'b	00011000,// -- a    **
8'b	00111100,// -- b   ****
8'b	00000000,// -- c
8'b	00000000,// -- d
8'b	00000000,// -- e
8'b	00000000},// -- f

{8'b	00000000,// -- 0 // O
8'b	00000000,// -- 1
8'b	01111100,// -- 2  *****
8'b	11000110,// -- 3 **   **
8'b	11000110,// -- 4 **   **
8'b	11000110,// -- 5 **   **
8'b	11000110,// -- 6 **   **
8'b	11000110,// -- 7 **   **
8'b	11000110,// -- 8 **   **
8'b	11000110,// -- 9 **   **
8'b	11000110,// -- a **   **
8'b	01111100,// -- b  *****
8'b	00000000,// -- c
8'b	00000000,// -- d
8'b	00000000,// -- e
8'b	00000000},// -- f

{8'b	00000000,// -- 0 // N
8'b	00000000,// -- 1
8'b	11000110,// -- 2 **   **
8'b	11100110,// -- 3 ***  **
8'b	11110110,// -- 4 **** **
8'b	11111110,// -- 5 *******
8'b	11011110,// -- 6 ** ****
8'b	11001110,// -- 7 **  ***
8'b	11000110,// -- 8 **   **
8'b	11000110,// -- 9 **   **
8'b	11000110,// -- a **   **
8'b	11000110,// -- b **   **
8'b	00000000,// -- c
8'b	00000000,// -- d
8'b	00000000,// -- e
8'b	00000000},// -- f

{8'b	00000000,// -- 0 // D
8'b	00000000,// -- 1
8'b	11111000,// -- 2 *****
8'b	01101100,// -- 3  ** **
8'b	01100110,// -- 4  **  **
8'b	01100110,// -- 5  **  **
8'b	01100110,// -- 6  **  **
8'b	01100110,// -- 7  **  **
8'b	01100110,// -- 8  **  **
8'b	01100110,// -- 9  **  **
8'b	01101100,// -- a  ** **
8'b	11111000,// -- b *****
8'b	00000000,// -- c
8'b	00000000,// -- d
8'b	00000000,// -- e
8'b	00000000},// -- f

{8'b	00000000,// -- 0 // M
8'b	00000000,// -- 1
8'b	11000011,// -- 2 **    **
8'b	11100111,// -- 3 ***  ***
8'b	11111111,// -- 4 ********
8'b	11111111,// -- 5 ********
8'b	11011011,// -- 6 ** ** **
8'b	11000011,// -- 7 **    **
8'b	11000011,// -- 8 **    **
8'b	11000011,// -- 9 **    **
8'b	11000011,// -- a **    **
8'b	11000011,// -- b **    **
8'b	00000000,// -- c
8'b	00000000,// -- d
8'b	00000000,// -- e
8'b	00000000},// -- f

{8'b	00000000,// -- 0 // I
8'b	00000000,// -- 1
8'b	00111100,// -- 2   ****
8'b	00011000,// -- 3    **
8'b	00011000,// -- 4    **
8'b	00011000,// -- 5    **
8'b	00011000,// -- 6    **
8'b	00011000,// -- 7    **
8'b	00011000,// -- 8    **
8'b	00011000,// -- 9    **
8'b	00011000,// -- a    **
8'b	00111100,// -- b   ****
8'b	00000000,// -- c
8'b	00000000,// -- d
8'b	00000000,// -- e
8'b	00000000},// -- f

{8'b	00000000,// -- 0 // Z
8'b	00000000,// -- 1
8'b	11111111,// -- 2 ********
8'b	11000011,// -- 3 **    **
8'b	10000110,// -- 4 *    **
8'b	00001100,// -- 5     **
8'b	00011000,// -- 6    **
8'b	00110000,// -- 7   **
8'b	01100000,// -- 8  **
8'b	11000001,// -- 9 **     *
8'b	11000011,// -- a **    **
8'b	11111111,// -- b ********
8'b	00000000,// -- c
8'b	00000000,// -- d
8'b	00000000,// -- e
8'b	00000000},// -- f

{8'b	00000000,// -- 0 // B
8'b	00000000,// -- 1
8'b	11111100,// -- 2 ******
8'b	01100110,// -- 3  **  **
8'b	01100110,// -- 4  **  **
8'b	01100110,// -- 5  **  **
8'b	01111100,// -- 6  *****
8'b	01100110,// -- 7  **  **
8'b	01100110,// -- 8  **  **
8'b	01100110,// -- 9  **  **
8'b	01100110,// -- a  **  **
8'b	11111100,// -- b ******
8'b	00000000,// -- c
8'b	00000000,// -- d
8'b	00000000,// -- e
8'b	00000000},// -- f

{8'b	00000000,// -- 0 // K
8'b	00000000,// -- 1
8'b	11100110,// -- 2 ***  **
8'b	01100110,// -- 3  **  **
8'b	01100110,// -- 4  **  **
8'b	01101100,// -- 5  ** **
8'b	01111000,// -- 6  ****
8'b	01111000,// -- 7  ****
8'b	01101100,// -- 8  ** **
8'b	01100110,// -- 9  **  **
8'b	01100110,// -- a  **  **
8'b	11100110,// -- b ***  **
8'b	00000000,// -- c
8'b	00000000,// -- d
8'b	00000000,// -- e
8'b	00000000},// -- f

{8'b	00000000,// -- 0 // Y
8'b	00000000,// -- 1
8'b	11000011,// -- 2 **    **
8'b	11000011,// -- 3 **    **
8'b	11000011,// -- 4 **    **
8'b	01100110,// -- 5  **  **
8'b	00111100,// -- 6   ****
8'b	00011000,// -- 7    **
8'b	00011000,// -- 8    **
8'b	00011000,// -- 9    **
8'b	00011000,// -- a    **
8'b	00111100,// -- b   ****
8'b	00000000,// -- c
8'b	00000000,// -- d
8'b	00000000,// -- e
8'b	00000000},// -- f

{8'b	00000000,// -- 0 // U
8'b	00000000,// -- 1
8'b	11000110,// -- 2 **   **
8'b	11000110,// -- 3 **   **
8'b	11000110,// -- 4 **   **
8'b	11000110,// -- 5 **   **
8'b	11000110,// -- 6 **   **
8'b	11000110,// -- 7 **   **
8'b	11000110,// -- 8 **   **
8'b	11000110,// -- 9 **   **
8'b	11000110,// -- a **   **
8'b	01111100,// -- b  *****
8'b	00000000,// -- c
8'b	00000000,// -- d
8'b	00000000,// -- e
8'b	00000000},// -- f

{8'b	00000000,// -- 0 // W
8'b	00000000,// -- 1
8'b	11000011,// -- 2 **    **
8'b	11000011,// -- 3 **    **
8'b	11000011,// -- 4 **    **
8'b	11000011,// -- 5 **    **
8'b	11000011,// -- 6 **    **
8'b	11011011,// -- 7 ** ** **
8'b	11011011,// -- 8 ** ** **
8'b	11111111,// -- 9 ********
8'b	01100110,// -- a  **  **
8'b	01100110,// -- b  **  **
8'b	00000000,// -- c
8'b	00000000,// -- d
8'b	00000000,// -- e
8'b	00000000},// -- f

{8'b	00000000,// -- 0 // L
8'b	00000000,// -- 1
8'b	11110000,// -- 2 ****
8'b	01100000,// -- 3  **
8'b	01100000,// -- 4  **
8'b	01100000,// -- 5  **
8'b	01100000,// -- 6  **
8'b	01100000,// -- 7  **
8'b	01100000,// -- 8  **
8'b	01100010,// -- 9  **   *
8'b	01100110,// -- a  **  **
8'b	11111110,// -- b *******
8'b	00000000,// -- c
8'b	00000000,// -- d
8'b	00000000,// -- e
8'b	00000000}// -- f
					
} ;				

// pipeline (ff) to get the pixel color from the array 	 

always_ff@(posedge clk or negedge resetN)
begin
	if(!resetN) begin
		drawingRequest <=	1'b0;
	end
	else begin
			drawingRequest <= (letter_bitmap[letter][offsetY/4][offsetX/4]) && (InsideRectangle == 1'b1 );	//get value from bitmap and enlarge ist size 4 times
	end 
end

assign RGBout = digit_color ; // this is a fixed color 

endmodule
